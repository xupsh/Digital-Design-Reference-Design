`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2014/10/30 22:27:12
// Design Name: 
// Module Name: BtoD
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module BtoD(
input[7:0]R_detect,G_detect,B_detect,
output reg[3:0]R_h,R_d,R_u,
output reg[3:0]G_h,G_d,G_u,
output reg[3:0]B_h,B_d,B_u
    );
 always@(*)begin
case (R_detect)
8'd0:begin R_h <=4'd0;R_d<=4'd0;R_u<=4'd0;end
8'd1:begin R_h <=4'd0;R_d<=4'd0;R_u<=4'd1;end
8'd2:begin R_h <=4'd0;R_d<=4'd0;R_u<=4'd2;end
8'd3:begin R_h <=4'd0;R_d<=4'd0;R_u<=4'd3;end
8'd4:begin R_h <=4'd0;R_d<=4'd0;R_u<=4'd4;end
8'd5:begin R_h <=4'd0;R_d<=4'd0;R_u<=4'd5;end
8'd6:begin R_h <=4'd0;R_d<=4'd0;R_u<=4'd6;end
8'd7:begin R_h <=4'd0;R_d<=4'd0;R_u<=4'd7;end
8'd8:begin R_h <=4'd0;R_d<=4'd0;R_u<=4'd8;end
8'd9:begin R_h <=4'd0;R_d<=4'd0;R_u<=4'd9;end
8'd10:begin R_h <=4'd0;R_d<=4'd1;R_u<=4'd0;end
8'd11:begin R_h <=4'd0;R_d<=4'd1;R_u<=4'd1;end
8'd12:begin R_h <=4'd0;R_d<=4'd1;R_u<=4'd2;end
8'd13:begin R_h <=4'd0;R_d<=4'd1;R_u<=4'd3;end
8'd14:begin R_h <=4'd0;R_d<=4'd1;R_u<=4'd4;end
8'd15:begin R_h <=4'd0;R_d<=4'd1;R_u<=4'd5;end
8'd16:begin R_h <=4'd0;R_d<=4'd1;R_u<=4'd6;end
8'd17:begin R_h <=4'd0;R_d<=4'd1;R_u<=4'd7;end
8'd18:begin R_h <=4'd0;R_d<=4'd1;R_u<=4'd8;end
8'd19:begin R_h <=4'd0;R_d<=4'd1;R_u<=4'd9;end
8'd20:begin R_h <=4'd0;R_d<=4'd2;R_u<=4'd0;end
8'd21:begin R_h <=4'd0;R_d<=4'd2;R_u<=4'd1;end
8'd22:begin R_h <=4'd0;R_d<=4'd2;R_u<=4'd2;end
8'd23:begin R_h <=4'd0;R_d<=4'd2;R_u<=4'd3;end
8'd24:begin R_h <=4'd0;R_d<=4'd2;R_u<=4'd4;end
8'd25:begin R_h <=4'd0;R_d<=4'd2;R_u<=4'd5;end
8'd26:begin R_h <=4'd0;R_d<=4'd2;R_u<=4'd6;end
8'd27:begin R_h <=4'd0;R_d<=4'd2;R_u<=4'd7;end
8'd28:begin R_h <=4'd0;R_d<=4'd2;R_u<=4'd8;end
8'd29:begin R_h <=4'd0;R_d<=4'd2;R_u<=4'd9;end
8'd30:begin R_h <=4'd0;R_d<=4'd3;R_u<=4'd0;end
8'd31:begin R_h <=4'd0;R_d<=4'd3;R_u<=4'd1;end
8'd32:begin R_h <=4'd0;R_d<=4'd3;R_u<=4'd2;end
8'd33:begin R_h <=4'd0;R_d<=4'd3;R_u<=4'd3;end
8'd34:begin R_h <=4'd0;R_d<=4'd3;R_u<=4'd4;end
8'd35:begin R_h <=4'd0;R_d<=4'd3;R_u<=4'd5;end
8'd36:begin R_h <=4'd0;R_d<=4'd3;R_u<=4'd6;end
8'd37:begin R_h <=4'd0;R_d<=4'd3;R_u<=4'd7;end
8'd38:begin R_h <=4'd0;R_d<=4'd3;R_u<=4'd8;end
8'd39:begin R_h <=4'd0;R_d<=4'd3;R_u<=4'd9;end
8'd40:begin R_h <=4'd0;R_d<=4'd4;R_u<=4'd0;end
8'd41:begin R_h <=4'd0;R_d<=4'd4;R_u<=4'd1;end
8'd42:begin R_h <=4'd0;R_d<=4'd4;R_u<=4'd2;end
8'd43:begin R_h <=4'd0;R_d<=4'd4;R_u<=4'd3;end
8'd44:begin R_h <=4'd0;R_d<=4'd4;R_u<=4'd4;end
8'd45:begin R_h <=4'd0;R_d<=4'd4;R_u<=4'd5;end
8'd46:begin R_h <=4'd0;R_d<=4'd4;R_u<=4'd6;end
8'd47:begin R_h <=4'd0;R_d<=4'd4;R_u<=4'd7;end
8'd48:begin R_h <=4'd0;R_d<=4'd4;R_u<=4'd8;end
8'd49:begin R_h <=4'd0;R_d<=4'd4;R_u<=4'd9;end
8'd50:begin R_h <=4'd0;R_d<=4'd5;R_u<=4'd0;end
8'd51:begin R_h <=4'd0;R_d<=4'd5;R_u<=4'd1;end
8'd52:begin R_h <=4'd0;R_d<=4'd5;R_u<=4'd2;end
8'd53:begin R_h <=4'd0;R_d<=4'd5;R_u<=4'd3;end
8'd54:begin R_h <=4'd0;R_d<=4'd5;R_u<=4'd4;end
8'd55:begin R_h <=4'd0;R_d<=4'd5;R_u<=4'd5;end
8'd56:begin R_h <=4'd0;R_d<=4'd5;R_u<=4'd6;end
8'd57:begin R_h <=4'd0;R_d<=4'd5;R_u<=4'd7;end
8'd58:begin R_h <=4'd0;R_d<=4'd5;R_u<=4'd8;end
8'd59:begin R_h <=4'd0;R_d<=4'd5;R_u<=4'd9;end
8'd60:begin R_h <=4'd0;R_d<=4'd6;R_u<=4'd0;end
8'd61:begin R_h <=4'd0;R_d<=4'd6;R_u<=4'd1;end
8'd62:begin R_h <=4'd0;R_d<=4'd6;R_u<=4'd2;end
8'd63:begin R_h <=4'd0;R_d<=4'd6;R_u<=4'd3;end
8'd64:begin R_h <=4'd0;R_d<=4'd6;R_u<=4'd4;end
8'd65:begin R_h <=4'd0;R_d<=4'd6;R_u<=4'd5;end
8'd66:begin R_h <=4'd0;R_d<=4'd6;R_u<=4'd6;end
8'd67:begin R_h <=4'd0;R_d<=4'd6;R_u<=4'd7;end
8'd68:begin R_h <=4'd0;R_d<=4'd6;R_u<=4'd8;end
8'd69:begin R_h <=4'd0;R_d<=4'd6;R_u<=4'd9;end
8'd70:begin R_h <=4'd0;R_d<=4'd7;R_u<=4'd0;end
8'd71:begin R_h <=4'd0;R_d<=4'd7;R_u<=4'd1;end
8'd72:begin R_h <=4'd0;R_d<=4'd7;R_u<=4'd2;end
8'd73:begin R_h <=4'd0;R_d<=4'd7;R_u<=4'd3;end
8'd74:begin R_h <=4'd0;R_d<=4'd7;R_u<=4'd4;end
8'd75:begin R_h <=4'd0;R_d<=4'd7;R_u<=4'd5;end
8'd76:begin R_h <=4'd0;R_d<=4'd7;R_u<=4'd6;end
8'd77:begin R_h <=4'd0;R_d<=4'd7;R_u<=4'd7;end
8'd78:begin R_h <=4'd0;R_d<=4'd7;R_u<=4'd8;end
8'd79:begin R_h <=4'd0;R_d<=4'd7;R_u<=4'd9;end
8'd80:begin R_h <=4'd0;R_d<=4'd8;R_u<=4'd0;end
8'd81:begin R_h <=4'd0;R_d<=4'd8;R_u<=4'd1;end
8'd82:begin R_h <=4'd0;R_d<=4'd8;R_u<=4'd2;end
8'd83:begin R_h <=4'd0;R_d<=4'd8;R_u<=4'd3;end
8'd84:begin R_h <=4'd0;R_d<=4'd8;R_u<=4'd4;end
8'd85:begin R_h <=4'd0;R_d<=4'd8;R_u<=4'd5;end
8'd86:begin R_h <=4'd0;R_d<=4'd8;R_u<=4'd6;end
8'd87:begin R_h <=4'd0;R_d<=4'd8;R_u<=4'd7;end
8'd88:begin R_h <=4'd0;R_d<=4'd8;R_u<=4'd8;end
8'd89:begin R_h <=4'd0;R_d<=4'd8;R_u<=4'd9;end
8'd90:begin R_h <=4'd0;R_d<=4'd9;R_u<=4'd0;end
8'd91:begin R_h <=4'd0;R_d<=4'd9;R_u<=4'd1;end
8'd92:begin R_h <=4'd0;R_d<=4'd9;R_u<=4'd2;end
8'd93:begin R_h <=4'd0;R_d<=4'd9;R_u<=4'd3;end
8'd94:begin R_h <=4'd0;R_d<=4'd9;R_u<=4'd4;end
8'd95:begin R_h <=4'd0;R_d<=4'd9;R_u<=4'd5;end
8'd96:begin R_h <=4'd0;R_d<=4'd9;R_u<=4'd6;end
8'd97:begin R_h <=4'd0;R_d<=4'd9;R_u<=4'd7;end
8'd98:begin R_h <=4'd0;R_d<=4'd9;R_u<=4'd8;end
8'd99:begin R_h <=4'd0;R_d<=4'd9;R_u<=4'd9;end
8'd100:begin R_h <=4'd1;R_d<=4'd0;R_u<=4'd0;end
8'd101:begin R_h <=4'd1;R_d<=4'd0;R_u<=4'd1;end
8'd102:begin R_h <=4'd1;R_d<=4'd0;R_u<=4'd2;end
8'd103:begin R_h <=4'd1;R_d<=4'd0;R_u<=4'd3;end
8'd104:begin R_h <=4'd1;R_d<=4'd0;R_u<=4'd4;end
8'd105:begin R_h <=4'd1;R_d<=4'd0;R_u<=4'd5;end
8'd106:begin R_h <=4'd1;R_d<=4'd0;R_u<=4'd6;end
8'd107:begin R_h <=4'd1;R_d<=4'd0;R_u<=4'd7;end
8'd108:begin R_h <=4'd1;R_d<=4'd0;R_u<=4'd8;end
8'd109:begin R_h <=4'd1;R_d<=4'd0;R_u<=4'd9;end
8'd110:begin R_h <=4'd1;R_d<=4'd1;R_u<=4'd0;end
8'd111:begin R_h <=4'd1;R_d<=4'd1;R_u<=4'd1;end
8'd112:begin R_h <=4'd1;R_d<=4'd1;R_u<=4'd2;end
8'd113:begin R_h <=4'd1;R_d<=4'd1;R_u<=4'd3;end
8'd114:begin R_h <=4'd1;R_d<=4'd1;R_u<=4'd4;end
8'd115:begin R_h <=4'd1;R_d<=4'd1;R_u<=4'd5;end
8'd116:begin R_h <=4'd1;R_d<=4'd1;R_u<=4'd6;end
8'd117:begin R_h <=4'd1;R_d<=4'd1;R_u<=4'd7;end
8'd118:begin R_h <=4'd1;R_d<=4'd1;R_u<=4'd8;end
8'd119:begin R_h <=4'd1;R_d<=4'd1;R_u<=4'd9;end
8'd120:begin R_h <=4'd1;R_d<=4'd2;R_u<=4'd0;end
8'd121:begin R_h <=4'd1;R_d<=4'd2;R_u<=4'd1;end
8'd122:begin R_h <=4'd1;R_d<=4'd2;R_u<=4'd2;end
8'd123:begin R_h <=4'd1;R_d<=4'd2;R_u<=4'd3;end
8'd124:begin R_h <=4'd1;R_d<=4'd2;R_u<=4'd4;end
8'd125:begin R_h <=4'd1;R_d<=4'd2;R_u<=4'd5;end
8'd126:begin R_h <=4'd1;R_d<=4'd2;R_u<=4'd6;end
8'd127:begin R_h <=4'd1;R_d<=4'd2;R_u<=4'd7;end
8'd128:begin R_h <=4'd1;R_d<=4'd2;R_u<=4'd8;end
8'd129:begin R_h <=4'd1;R_d<=4'd2;R_u<=4'd9;end
8'd130:begin R_h <=4'd1;R_d<=4'd3;R_u<=4'd0;end
8'd131:begin R_h <=4'd1;R_d<=4'd3;R_u<=4'd1;end
8'd132:begin R_h <=4'd1;R_d<=4'd3;R_u<=4'd2;end
8'd133:begin R_h <=4'd1;R_d<=4'd3;R_u<=4'd3;end
8'd134:begin R_h <=4'd1;R_d<=4'd3;R_u<=4'd4;end
8'd135:begin R_h <=4'd1;R_d<=4'd3;R_u<=4'd5;end
8'd136:begin R_h <=4'd1;R_d<=4'd3;R_u<=4'd6;end
8'd137:begin R_h <=4'd1;R_d<=4'd3;R_u<=4'd7;end
8'd138:begin R_h <=4'd1;R_d<=4'd3;R_u<=4'd8;end
8'd139:begin R_h <=4'd1;R_d<=4'd3;R_u<=4'd9;end
8'd140:begin R_h <=4'd1;R_d<=4'd4;R_u<=4'd0;end
8'd141:begin R_h <=4'd1;R_d<=4'd4;R_u<=4'd1;end
8'd142:begin R_h <=4'd1;R_d<=4'd4;R_u<=4'd2;end
8'd143:begin R_h <=4'd1;R_d<=4'd4;R_u<=4'd3;end
8'd144:begin R_h <=4'd1;R_d<=4'd4;R_u<=4'd4;end
8'd145:begin R_h <=4'd1;R_d<=4'd4;R_u<=4'd5;end
8'd146:begin R_h <=4'd1;R_d<=4'd4;R_u<=4'd6;end
8'd147:begin R_h <=4'd1;R_d<=4'd4;R_u<=4'd7;end
8'd148:begin R_h <=4'd1;R_d<=4'd4;R_u<=4'd8;end
8'd149:begin R_h <=4'd1;R_d<=4'd4;R_u<=4'd9;end
8'd150:begin R_h <=4'd1;R_d<=4'd5;R_u<=4'd0;end
8'd151:begin R_h <=4'd1;R_d<=4'd5;R_u<=4'd1;end
8'd152:begin R_h <=4'd1;R_d<=4'd5;R_u<=4'd2;end
8'd153:begin R_h <=4'd1;R_d<=4'd5;R_u<=4'd3;end
8'd154:begin R_h <=4'd1;R_d<=4'd5;R_u<=4'd4;end
8'd155:begin R_h <=4'd1;R_d<=4'd5;R_u<=4'd5;end
8'd156:begin R_h <=4'd1;R_d<=4'd5;R_u<=4'd6;end
8'd157:begin R_h <=4'd1;R_d<=4'd5;R_u<=4'd7;end
8'd158:begin R_h <=4'd1;R_d<=4'd5;R_u<=4'd8;end
8'd159:begin R_h <=4'd1;R_d<=4'd5;R_u<=4'd9;end
8'd160:begin R_h <=4'd1;R_d<=4'd6;R_u<=4'd0;end
8'd161:begin R_h <=4'd1;R_d<=4'd6;R_u<=4'd1;end
8'd162:begin R_h <=4'd1;R_d<=4'd6;R_u<=4'd2;end
8'd163:begin R_h <=4'd1;R_d<=4'd6;R_u<=4'd3;end
8'd164:begin R_h <=4'd1;R_d<=4'd6;R_u<=4'd4;end
8'd165:begin R_h <=4'd1;R_d<=4'd6;R_u<=4'd5;end
8'd166:begin R_h <=4'd1;R_d<=4'd6;R_u<=4'd6;end
8'd167:begin R_h <=4'd1;R_d<=4'd6;R_u<=4'd7;end
8'd168:begin R_h <=4'd1;R_d<=4'd6;R_u<=4'd8;end
8'd169:begin R_h <=4'd1;R_d<=4'd6;R_u<=4'd9;end
8'd170:begin R_h <=4'd1;R_d<=4'd7;R_u<=4'd0;end
8'd171:begin R_h <=4'd1;R_d<=4'd7;R_u<=4'd1;end
8'd172:begin R_h <=4'd1;R_d<=4'd7;R_u<=4'd2;end
8'd173:begin R_h <=4'd1;R_d<=4'd7;R_u<=4'd3;end
8'd174:begin R_h <=4'd1;R_d<=4'd7;R_u<=4'd4;end
8'd175:begin R_h <=4'd1;R_d<=4'd7;R_u<=4'd5;end
8'd176:begin R_h <=4'd1;R_d<=4'd7;R_u<=4'd6;end
8'd177:begin R_h <=4'd1;R_d<=4'd7;R_u<=4'd7;end
8'd178:begin R_h <=4'd1;R_d<=4'd7;R_u<=4'd8;end
8'd179:begin R_h <=4'd1;R_d<=4'd7;R_u<=4'd9;end
8'd180:begin R_h <=4'd1;R_d<=4'd8;R_u<=4'd0;end
8'd181:begin R_h <=4'd1;R_d<=4'd8;R_u<=4'd1;end
8'd182:begin R_h <=4'd1;R_d<=4'd8;R_u<=4'd2;end
8'd183:begin R_h <=4'd1;R_d<=4'd8;R_u<=4'd3;end
8'd184:begin R_h <=4'd1;R_d<=4'd8;R_u<=4'd4;end
8'd185:begin R_h <=4'd1;R_d<=4'd8;R_u<=4'd5;end
8'd186:begin R_h <=4'd1;R_d<=4'd8;R_u<=4'd6;end
8'd187:begin R_h <=4'd1;R_d<=4'd8;R_u<=4'd7;end
8'd188:begin R_h <=4'd1;R_d<=4'd8;R_u<=4'd8;end
8'd189:begin R_h <=4'd1;R_d<=4'd8;R_u<=4'd9;end
8'd190:begin R_h <=4'd1;R_d<=4'd9;R_u<=4'd0;end
8'd191:begin R_h <=4'd1;R_d<=4'd9;R_u<=4'd1;end
8'd192:begin R_h <=4'd1;R_d<=4'd9;R_u<=4'd2;end
8'd193:begin R_h <=4'd1;R_d<=4'd9;R_u<=4'd3;end
8'd194:begin R_h <=4'd1;R_d<=4'd9;R_u<=4'd4;end
8'd195:begin R_h <=4'd1;R_d<=4'd9;R_u<=4'd5;end
8'd196:begin R_h <=4'd1;R_d<=4'd9;R_u<=4'd6;end
8'd197:begin R_h <=4'd1;R_d<=4'd9;R_u<=4'd7;end
8'd198:begin R_h <=4'd1;R_d<=4'd9;R_u<=4'd8;end
8'd199:begin R_h <=4'd1;R_d<=4'd9;R_u<=4'd9;end
8'd200:begin R_h <=4'd2;R_d<=4'd0;R_u<=4'd0;end
8'd201:begin R_h <=4'd2;R_d<=4'd0;R_u<=4'd1;end
8'd202:begin R_h <=4'd2;R_d<=4'd0;R_u<=4'd2;end
8'd203:begin R_h <=4'd2;R_d<=4'd0;R_u<=4'd3;end
8'd204:begin R_h <=4'd2;R_d<=4'd0;R_u<=4'd4;end
8'd205:begin R_h <=4'd2;R_d<=4'd0;R_u<=4'd5;end
8'd206:begin R_h <=4'd2;R_d<=4'd0;R_u<=4'd6;end
8'd207:begin R_h <=4'd2;R_d<=4'd0;R_u<=4'd7;end
8'd208:begin R_h <=4'd2;R_d<=4'd0;R_u<=4'd8;end
8'd209:begin R_h <=4'd2;R_d<=4'd0;R_u<=4'd9;end
8'd210:begin R_h <=4'd2;R_d<=4'd1;R_u<=4'd0;end
8'd211:begin R_h <=4'd2;R_d<=4'd1;R_u<=4'd1;end
8'd212:begin R_h <=4'd2;R_d<=4'd1;R_u<=4'd2;end
8'd213:begin R_h <=4'd2;R_d<=4'd1;R_u<=4'd3;end
8'd214:begin R_h <=4'd2;R_d<=4'd1;R_u<=4'd4;end
8'd215:begin R_h <=4'd2;R_d<=4'd1;R_u<=4'd5;end
8'd216:begin R_h <=4'd2;R_d<=4'd1;R_u<=4'd6;end
8'd217:begin R_h <=4'd2;R_d<=4'd1;R_u<=4'd7;end
8'd218:begin R_h <=4'd2;R_d<=4'd1;R_u<=4'd8;end
8'd219:begin R_h <=4'd2;R_d<=4'd1;R_u<=4'd9;end
8'd220:begin R_h <=4'd2;R_d<=4'd2;R_u<=4'd0;end
8'd221:begin R_h <=4'd2;R_d<=4'd2;R_u<=4'd1;end
8'd222:begin R_h <=4'd2;R_d<=4'd2;R_u<=4'd2;end
8'd223:begin R_h <=4'd2;R_d<=4'd2;R_u<=4'd3;end
8'd224:begin R_h <=4'd2;R_d<=4'd2;R_u<=4'd4;end
8'd225:begin R_h <=4'd2;R_d<=4'd2;R_u<=4'd5;end
8'd226:begin R_h <=4'd2;R_d<=4'd2;R_u<=4'd6;end
8'd227:begin R_h <=4'd2;R_d<=4'd2;R_u<=4'd7;end
8'd228:begin R_h <=4'd2;R_d<=4'd2;R_u<=4'd8;end
8'd229:begin R_h <=4'd2;R_d<=4'd2;R_u<=4'd9;end
8'd230:begin R_h <=4'd2;R_d<=4'd3;R_u<=4'd0;end
8'd231:begin R_h <=4'd2;R_d<=4'd3;R_u<=4'd1;end
8'd232:begin R_h <=4'd2;R_d<=4'd3;R_u<=4'd2;end
8'd233:begin R_h <=4'd2;R_d<=4'd3;R_u<=4'd3;end
8'd234:begin R_h <=4'd2;R_d<=4'd3;R_u<=4'd4;end
8'd235:begin R_h <=4'd2;R_d<=4'd3;R_u<=4'd5;end
8'd236:begin R_h <=4'd2;R_d<=4'd3;R_u<=4'd6;end
8'd237:begin R_h <=4'd2;R_d<=4'd3;R_u<=4'd7;end
8'd238:begin R_h <=4'd2;R_d<=4'd3;R_u<=4'd8;end
8'd239:begin R_h <=4'd2;R_d<=4'd3;R_u<=4'd9;end
8'd240:begin R_h <=4'd2;R_d<=4'd4;R_u<=4'd0;end
8'd241:begin R_h <=4'd2;R_d<=4'd4;R_u<=4'd1;end
8'd242:begin R_h <=4'd2;R_d<=4'd4;R_u<=4'd2;end
8'd243:begin R_h <=4'd2;R_d<=4'd4;R_u<=4'd3;end
8'd244:begin R_h <=4'd2;R_d<=4'd4;R_u<=4'd4;end
8'd245:begin R_h <=4'd2;R_d<=4'd4;R_u<=4'd5;end
8'd246:begin R_h <=4'd2;R_d<=4'd4;R_u<=4'd6;end
8'd247:begin R_h <=4'd2;R_d<=4'd4;R_u<=4'd7;end
8'd248:begin R_h <=4'd2;R_d<=4'd4;R_u<=4'd8;end
8'd249:begin R_h <=4'd2;R_d<=4'd4;R_u<=4'd9;end
8'd250:begin R_h <=4'd2;R_d<=4'd5;R_u<=4'd0;end
8'd251:begin R_h <=4'd2;R_d<=4'd5;R_u<=4'd1;end
8'd252:begin R_h <=4'd2;R_d<=4'd5;R_u<=4'd2;end
8'd253:begin R_h <=4'd2;R_d<=4'd5;R_u<=4'd3;end
8'd254:begin R_h <=4'd2;R_d<=4'd5;R_u<=4'd4;end
8'd255:begin R_h <=4'd2;R_d<=4'd5;R_u<=4'd5;end
endcase
end

always@(*)begin
case (G_detect)
8'd0:begin G_h <=4'd0;G_d<=4'd0;G_u<=4'd0;end
8'd1:begin G_h <=4'd0;G_d<=4'd0;G_u<=4'd1;end
8'd2:begin G_h <=4'd0;G_d<=4'd0;G_u<=4'd2;end
8'd3:begin G_h <=4'd0;G_d<=4'd0;G_u<=4'd3;end
8'd4:begin G_h <=4'd0;G_d<=4'd0;G_u<=4'd4;end
8'd5:begin G_h <=4'd0;G_d<=4'd0;G_u<=4'd5;end
8'd6:begin G_h <=4'd0;G_d<=4'd0;G_u<=4'd6;end
8'd7:begin G_h <=4'd0;G_d<=4'd0;G_u<=4'd7;end
8'd8:begin G_h <=4'd0;G_d<=4'd0;G_u<=4'd8;end
8'd9:begin G_h <=4'd0;G_d<=4'd0;G_u<=4'd9;end
8'd10:begin G_h <=4'd0;G_d<=4'd1;G_u<=4'd0;end
8'd11:begin G_h <=4'd0;G_d<=4'd1;G_u<=4'd1;end
8'd12:begin G_h <=4'd0;G_d<=4'd1;G_u<=4'd2;end
8'd13:begin G_h <=4'd0;G_d<=4'd1;G_u<=4'd3;end
8'd14:begin G_h <=4'd0;G_d<=4'd1;G_u<=4'd4;end
8'd15:begin G_h <=4'd0;G_d<=4'd1;G_u<=4'd5;end
8'd16:begin G_h <=4'd0;G_d<=4'd1;G_u<=4'd6;end
8'd17:begin G_h <=4'd0;G_d<=4'd1;G_u<=4'd7;end
8'd18:begin G_h <=4'd0;G_d<=4'd1;G_u<=4'd8;end
8'd19:begin G_h <=4'd0;G_d<=4'd1;G_u<=4'd9;end
8'd20:begin G_h <=4'd0;G_d<=4'd2;G_u<=4'd0;end
8'd21:begin G_h <=4'd0;G_d<=4'd2;G_u<=4'd1;end
8'd22:begin G_h <=4'd0;G_d<=4'd2;G_u<=4'd2;end
8'd23:begin G_h <=4'd0;G_d<=4'd2;G_u<=4'd3;end
8'd24:begin G_h <=4'd0;G_d<=4'd2;G_u<=4'd4;end
8'd25:begin G_h <=4'd0;G_d<=4'd2;G_u<=4'd5;end
8'd26:begin G_h <=4'd0;G_d<=4'd2;G_u<=4'd6;end
8'd27:begin G_h <=4'd0;G_d<=4'd2;G_u<=4'd7;end
8'd28:begin G_h <=4'd0;G_d<=4'd2;G_u<=4'd8;end
8'd29:begin G_h <=4'd0;G_d<=4'd2;G_u<=4'd9;end
8'd30:begin G_h <=4'd0;G_d<=4'd3;G_u<=4'd0;end
8'd31:begin G_h <=4'd0;G_d<=4'd3;G_u<=4'd1;end
8'd32:begin G_h <=4'd0;G_d<=4'd3;G_u<=4'd2;end
8'd33:begin G_h <=4'd0;G_d<=4'd3;G_u<=4'd3;end
8'd34:begin G_h <=4'd0;G_d<=4'd3;G_u<=4'd4;end
8'd35:begin G_h <=4'd0;G_d<=4'd3;G_u<=4'd5;end
8'd36:begin G_h <=4'd0;G_d<=4'd3;G_u<=4'd6;end
8'd37:begin G_h <=4'd0;G_d<=4'd3;G_u<=4'd7;end
8'd38:begin G_h <=4'd0;G_d<=4'd3;G_u<=4'd8;end
8'd39:begin G_h <=4'd0;G_d<=4'd3;G_u<=4'd9;end
8'd40:begin G_h <=4'd0;G_d<=4'd4;G_u<=4'd0;end
8'd41:begin G_h <=4'd0;G_d<=4'd4;G_u<=4'd1;end
8'd42:begin G_h <=4'd0;G_d<=4'd4;G_u<=4'd2;end
8'd43:begin G_h <=4'd0;G_d<=4'd4;G_u<=4'd3;end
8'd44:begin G_h <=4'd0;G_d<=4'd4;G_u<=4'd4;end
8'd45:begin G_h <=4'd0;G_d<=4'd4;G_u<=4'd5;end
8'd46:begin G_h <=4'd0;G_d<=4'd4;G_u<=4'd6;end
8'd47:begin G_h <=4'd0;G_d<=4'd4;G_u<=4'd7;end
8'd48:begin G_h <=4'd0;G_d<=4'd4;G_u<=4'd8;end
8'd49:begin G_h <=4'd0;G_d<=4'd4;G_u<=4'd9;end
8'd50:begin G_h <=4'd0;G_d<=4'd5;G_u<=4'd0;end
8'd51:begin G_h <=4'd0;G_d<=4'd5;G_u<=4'd1;end
8'd52:begin G_h <=4'd0;G_d<=4'd5;G_u<=4'd2;end
8'd53:begin G_h <=4'd0;G_d<=4'd5;G_u<=4'd3;end
8'd54:begin G_h <=4'd0;G_d<=4'd5;G_u<=4'd4;end
8'd55:begin G_h <=4'd0;G_d<=4'd5;G_u<=4'd5;end
8'd56:begin G_h <=4'd0;G_d<=4'd5;G_u<=4'd6;end
8'd57:begin G_h <=4'd0;G_d<=4'd5;G_u<=4'd7;end
8'd58:begin G_h <=4'd0;G_d<=4'd5;G_u<=4'd8;end
8'd59:begin G_h <=4'd0;G_d<=4'd5;G_u<=4'd9;end
8'd60:begin G_h <=4'd0;G_d<=4'd6;G_u<=4'd0;end
8'd61:begin G_h <=4'd0;G_d<=4'd6;G_u<=4'd1;end
8'd62:begin G_h <=4'd0;G_d<=4'd6;G_u<=4'd2;end
8'd63:begin G_h <=4'd0;G_d<=4'd6;G_u<=4'd3;end
8'd64:begin G_h <=4'd0;G_d<=4'd6;G_u<=4'd4;end
8'd65:begin G_h <=4'd0;G_d<=4'd6;G_u<=4'd5;end
8'd66:begin G_h <=4'd0;G_d<=4'd6;G_u<=4'd6;end
8'd67:begin G_h <=4'd0;G_d<=4'd6;G_u<=4'd7;end
8'd68:begin G_h <=4'd0;G_d<=4'd6;G_u<=4'd8;end
8'd69:begin G_h <=4'd0;G_d<=4'd6;G_u<=4'd9;end
8'd70:begin G_h <=4'd0;G_d<=4'd7;G_u<=4'd0;end
8'd71:begin G_h <=4'd0;G_d<=4'd7;G_u<=4'd1;end
8'd72:begin G_h <=4'd0;G_d<=4'd7;G_u<=4'd2;end
8'd73:begin G_h <=4'd0;G_d<=4'd7;G_u<=4'd3;end
8'd74:begin G_h <=4'd0;G_d<=4'd7;G_u<=4'd4;end
8'd75:begin G_h <=4'd0;G_d<=4'd7;G_u<=4'd5;end
8'd76:begin G_h <=4'd0;G_d<=4'd7;G_u<=4'd6;end
8'd77:begin G_h <=4'd0;G_d<=4'd7;G_u<=4'd7;end
8'd78:begin G_h <=4'd0;G_d<=4'd7;G_u<=4'd8;end
8'd79:begin G_h <=4'd0;G_d<=4'd7;G_u<=4'd9;end
8'd80:begin G_h <=4'd0;G_d<=4'd8;G_u<=4'd0;end
8'd81:begin G_h <=4'd0;G_d<=4'd8;G_u<=4'd1;end
8'd82:begin G_h <=4'd0;G_d<=4'd8;G_u<=4'd2;end
8'd83:begin G_h <=4'd0;G_d<=4'd8;G_u<=4'd3;end
8'd84:begin G_h <=4'd0;G_d<=4'd8;G_u<=4'd4;end
8'd85:begin G_h <=4'd0;G_d<=4'd8;G_u<=4'd5;end
8'd86:begin G_h <=4'd0;G_d<=4'd8;G_u<=4'd6;end
8'd87:begin G_h <=4'd0;G_d<=4'd8;G_u<=4'd7;end
8'd88:begin G_h <=4'd0;G_d<=4'd8;G_u<=4'd8;end
8'd89:begin G_h <=4'd0;G_d<=4'd8;G_u<=4'd9;end
8'd90:begin G_h <=4'd0;G_d<=4'd9;G_u<=4'd0;end
8'd91:begin G_h <=4'd0;G_d<=4'd9;G_u<=4'd1;end
8'd92:begin G_h <=4'd0;G_d<=4'd9;G_u<=4'd2;end
8'd93:begin G_h <=4'd0;G_d<=4'd9;G_u<=4'd3;end
8'd94:begin G_h <=4'd0;G_d<=4'd9;G_u<=4'd4;end
8'd95:begin G_h <=4'd0;G_d<=4'd9;G_u<=4'd5;end
8'd96:begin G_h <=4'd0;G_d<=4'd9;G_u<=4'd6;end
8'd97:begin G_h <=4'd0;G_d<=4'd9;G_u<=4'd7;end
8'd98:begin G_h <=4'd0;G_d<=4'd9;G_u<=4'd8;end
8'd99:begin G_h <=4'd0;G_d<=4'd9;G_u<=4'd9;end
8'd100:begin G_h <=4'd1;G_d<=4'd0;G_u<=4'd0;end
8'd101:begin G_h <=4'd1;G_d<=4'd0;G_u<=4'd1;end
8'd102:begin G_h <=4'd1;G_d<=4'd0;G_u<=4'd2;end
8'd103:begin G_h <=4'd1;G_d<=4'd0;G_u<=4'd3;end
8'd104:begin G_h <=4'd1;G_d<=4'd0;G_u<=4'd4;end
8'd105:begin G_h <=4'd1;G_d<=4'd0;G_u<=4'd5;end
8'd106:begin G_h <=4'd1;G_d<=4'd0;G_u<=4'd6;end
8'd107:begin G_h <=4'd1;G_d<=4'd0;G_u<=4'd7;end
8'd108:begin G_h <=4'd1;G_d<=4'd0;G_u<=4'd8;end
8'd109:begin G_h <=4'd1;G_d<=4'd0;G_u<=4'd9;end
8'd110:begin G_h <=4'd1;G_d<=4'd1;G_u<=4'd0;end
8'd111:begin G_h <=4'd1;G_d<=4'd1;G_u<=4'd1;end
8'd112:begin G_h <=4'd1;G_d<=4'd1;G_u<=4'd2;end
8'd113:begin G_h <=4'd1;G_d<=4'd1;G_u<=4'd3;end
8'd114:begin G_h <=4'd1;G_d<=4'd1;G_u<=4'd4;end
8'd115:begin G_h <=4'd1;G_d<=4'd1;G_u<=4'd5;end
8'd116:begin G_h <=4'd1;G_d<=4'd1;G_u<=4'd6;end
8'd117:begin G_h <=4'd1;G_d<=4'd1;G_u<=4'd7;end
8'd118:begin G_h <=4'd1;G_d<=4'd1;G_u<=4'd8;end
8'd119:begin G_h <=4'd1;G_d<=4'd1;G_u<=4'd9;end
8'd120:begin G_h <=4'd1;G_d<=4'd2;G_u<=4'd0;end
8'd121:begin G_h <=4'd1;G_d<=4'd2;G_u<=4'd1;end
8'd122:begin G_h <=4'd1;G_d<=4'd2;G_u<=4'd2;end
8'd123:begin G_h <=4'd1;G_d<=4'd2;G_u<=4'd3;end
8'd124:begin G_h <=4'd1;G_d<=4'd2;G_u<=4'd4;end
8'd125:begin G_h <=4'd1;G_d<=4'd2;G_u<=4'd5;end
8'd126:begin G_h <=4'd1;G_d<=4'd2;G_u<=4'd6;end
8'd127:begin G_h <=4'd1;G_d<=4'd2;G_u<=4'd7;end
8'd128:begin G_h <=4'd1;G_d<=4'd2;G_u<=4'd8;end
8'd129:begin G_h <=4'd1;G_d<=4'd2;G_u<=4'd9;end
8'd130:begin G_h <=4'd1;G_d<=4'd3;G_u<=4'd0;end
8'd131:begin G_h <=4'd1;G_d<=4'd3;G_u<=4'd1;end
8'd132:begin G_h <=4'd1;G_d<=4'd3;G_u<=4'd2;end
8'd133:begin G_h <=4'd1;G_d<=4'd3;G_u<=4'd3;end
8'd134:begin G_h <=4'd1;G_d<=4'd3;G_u<=4'd4;end
8'd135:begin G_h <=4'd1;G_d<=4'd3;G_u<=4'd5;end
8'd136:begin G_h <=4'd1;G_d<=4'd3;G_u<=4'd6;end
8'd137:begin G_h <=4'd1;G_d<=4'd3;G_u<=4'd7;end
8'd138:begin G_h <=4'd1;G_d<=4'd3;G_u<=4'd8;end
8'd139:begin G_h <=4'd1;G_d<=4'd3;G_u<=4'd9;end
8'd140:begin G_h <=4'd1;G_d<=4'd4;G_u<=4'd0;end
8'd141:begin G_h <=4'd1;G_d<=4'd4;G_u<=4'd1;end
8'd142:begin G_h <=4'd1;G_d<=4'd4;G_u<=4'd2;end
8'd143:begin G_h <=4'd1;G_d<=4'd4;G_u<=4'd3;end
8'd144:begin G_h <=4'd1;G_d<=4'd4;G_u<=4'd4;end
8'd145:begin G_h <=4'd1;G_d<=4'd4;G_u<=4'd5;end
8'd146:begin G_h <=4'd1;G_d<=4'd4;G_u<=4'd6;end
8'd147:begin G_h <=4'd1;G_d<=4'd4;G_u<=4'd7;end
8'd148:begin G_h <=4'd1;G_d<=4'd4;G_u<=4'd8;end
8'd149:begin G_h <=4'd1;G_d<=4'd4;G_u<=4'd9;end
8'd150:begin G_h <=4'd1;G_d<=4'd5;G_u<=4'd0;end
8'd151:begin G_h <=4'd1;G_d<=4'd5;G_u<=4'd1;end
8'd152:begin G_h <=4'd1;G_d<=4'd5;G_u<=4'd2;end
8'd153:begin G_h <=4'd1;G_d<=4'd5;G_u<=4'd3;end
8'd154:begin G_h <=4'd1;G_d<=4'd5;G_u<=4'd4;end
8'd155:begin G_h <=4'd1;G_d<=4'd5;G_u<=4'd5;end
8'd156:begin G_h <=4'd1;G_d<=4'd5;G_u<=4'd6;end
8'd157:begin G_h <=4'd1;G_d<=4'd5;G_u<=4'd7;end
8'd158:begin G_h <=4'd1;G_d<=4'd5;G_u<=4'd8;end
8'd159:begin G_h <=4'd1;G_d<=4'd5;G_u<=4'd9;end
8'd160:begin G_h <=4'd1;G_d<=4'd6;G_u<=4'd0;end
8'd161:begin G_h <=4'd1;G_d<=4'd6;G_u<=4'd1;end
8'd162:begin G_h <=4'd1;G_d<=4'd6;G_u<=4'd2;end
8'd163:begin G_h <=4'd1;G_d<=4'd6;G_u<=4'd3;end
8'd164:begin G_h <=4'd1;G_d<=4'd6;G_u<=4'd4;end
8'd165:begin G_h <=4'd1;G_d<=4'd6;G_u<=4'd5;end
8'd166:begin G_h <=4'd1;G_d<=4'd6;G_u<=4'd6;end
8'd167:begin G_h <=4'd1;G_d<=4'd6;G_u<=4'd7;end
8'd168:begin G_h <=4'd1;G_d<=4'd6;G_u<=4'd8;end
8'd169:begin G_h <=4'd1;G_d<=4'd6;G_u<=4'd9;end
8'd170:begin G_h <=4'd1;G_d<=4'd7;G_u<=4'd0;end
8'd171:begin G_h <=4'd1;G_d<=4'd7;G_u<=4'd1;end
8'd172:begin G_h <=4'd1;G_d<=4'd7;G_u<=4'd2;end
8'd173:begin G_h <=4'd1;G_d<=4'd7;G_u<=4'd3;end
8'd174:begin G_h <=4'd1;G_d<=4'd7;G_u<=4'd4;end
8'd175:begin G_h <=4'd1;G_d<=4'd7;G_u<=4'd5;end
8'd176:begin G_h <=4'd1;G_d<=4'd7;G_u<=4'd6;end
8'd177:begin G_h <=4'd1;G_d<=4'd7;G_u<=4'd7;end
8'd178:begin G_h <=4'd1;G_d<=4'd7;G_u<=4'd8;end
8'd179:begin G_h <=4'd1;G_d<=4'd7;G_u<=4'd9;end
8'd180:begin G_h <=4'd1;G_d<=4'd8;G_u<=4'd0;end
8'd181:begin G_h <=4'd1;G_d<=4'd8;G_u<=4'd1;end
8'd182:begin G_h <=4'd1;G_d<=4'd8;G_u<=4'd2;end
8'd183:begin G_h <=4'd1;G_d<=4'd8;G_u<=4'd3;end
8'd184:begin G_h <=4'd1;G_d<=4'd8;G_u<=4'd4;end
8'd185:begin G_h <=4'd1;G_d<=4'd8;G_u<=4'd5;end
8'd186:begin G_h <=4'd1;G_d<=4'd8;G_u<=4'd6;end
8'd187:begin G_h <=4'd1;G_d<=4'd8;G_u<=4'd7;end
8'd188:begin G_h <=4'd1;G_d<=4'd8;G_u<=4'd8;end
8'd189:begin G_h <=4'd1;G_d<=4'd8;G_u<=4'd9;end
8'd190:begin G_h <=4'd1;G_d<=4'd9;G_u<=4'd0;end
8'd191:begin G_h <=4'd1;G_d<=4'd9;G_u<=4'd1;end
8'd192:begin G_h <=4'd1;G_d<=4'd9;G_u<=4'd2;end
8'd193:begin G_h <=4'd1;G_d<=4'd9;G_u<=4'd3;end
8'd194:begin G_h <=4'd1;G_d<=4'd9;G_u<=4'd4;end
8'd195:begin G_h <=4'd1;G_d<=4'd9;G_u<=4'd5;end
8'd196:begin G_h <=4'd1;G_d<=4'd9;G_u<=4'd6;end
8'd197:begin G_h <=4'd1;G_d<=4'd9;G_u<=4'd7;end
8'd198:begin G_h <=4'd1;G_d<=4'd9;G_u<=4'd8;end
8'd199:begin G_h <=4'd1;G_d<=4'd9;G_u<=4'd9;end
8'd200:begin G_h <=4'd2;G_d<=4'd0;G_u<=4'd0;end
8'd201:begin G_h <=4'd2;G_d<=4'd0;G_u<=4'd1;end
8'd202:begin G_h <=4'd2;G_d<=4'd0;G_u<=4'd2;end
8'd203:begin G_h <=4'd2;G_d<=4'd0;G_u<=4'd3;end
8'd204:begin G_h <=4'd2;G_d<=4'd0;G_u<=4'd4;end
8'd205:begin G_h <=4'd2;G_d<=4'd0;G_u<=4'd5;end
8'd206:begin G_h <=4'd2;G_d<=4'd0;G_u<=4'd6;end
8'd207:begin G_h <=4'd2;G_d<=4'd0;G_u<=4'd7;end
8'd208:begin G_h <=4'd2;G_d<=4'd0;G_u<=4'd8;end
8'd209:begin G_h <=4'd2;G_d<=4'd0;G_u<=4'd9;end
8'd210:begin G_h <=4'd2;G_d<=4'd1;G_u<=4'd0;end
8'd211:begin G_h <=4'd2;G_d<=4'd1;G_u<=4'd1;end
8'd212:begin G_h <=4'd2;G_d<=4'd1;G_u<=4'd2;end
8'd213:begin G_h <=4'd2;G_d<=4'd1;G_u<=4'd3;end
8'd214:begin G_h <=4'd2;G_d<=4'd1;G_u<=4'd4;end
8'd215:begin G_h <=4'd2;G_d<=4'd1;G_u<=4'd5;end
8'd216:begin G_h <=4'd2;G_d<=4'd1;G_u<=4'd6;end
8'd217:begin G_h <=4'd2;G_d<=4'd1;G_u<=4'd7;end
8'd218:begin G_h <=4'd2;G_d<=4'd1;G_u<=4'd8;end
8'd219:begin G_h <=4'd2;G_d<=4'd1;G_u<=4'd9;end
8'd220:begin G_h <=4'd2;G_d<=4'd2;G_u<=4'd0;end
8'd221:begin G_h <=4'd2;G_d<=4'd2;G_u<=4'd1;end
8'd222:begin G_h <=4'd2;G_d<=4'd2;G_u<=4'd2;end
8'd223:begin G_h <=4'd2;G_d<=4'd2;G_u<=4'd3;end
8'd224:begin G_h <=4'd2;G_d<=4'd2;G_u<=4'd4;end
8'd225:begin G_h <=4'd2;G_d<=4'd2;G_u<=4'd5;end
8'd226:begin G_h <=4'd2;G_d<=4'd2;G_u<=4'd6;end
8'd227:begin G_h <=4'd2;G_d<=4'd2;G_u<=4'd7;end
8'd228:begin G_h <=4'd2;G_d<=4'd2;G_u<=4'd8;end
8'd229:begin G_h <=4'd2;G_d<=4'd2;G_u<=4'd9;end
8'd230:begin G_h <=4'd2;G_d<=4'd3;G_u<=4'd0;end
8'd231:begin G_h <=4'd2;G_d<=4'd3;G_u<=4'd1;end
8'd232:begin G_h <=4'd2;G_d<=4'd3;G_u<=4'd2;end
8'd233:begin G_h <=4'd2;G_d<=4'd3;G_u<=4'd3;end
8'd234:begin G_h <=4'd2;G_d<=4'd3;G_u<=4'd4;end
8'd235:begin G_h <=4'd2;G_d<=4'd3;G_u<=4'd5;end
8'd236:begin G_h <=4'd2;G_d<=4'd3;G_u<=4'd6;end
8'd237:begin G_h <=4'd2;G_d<=4'd3;G_u<=4'd7;end
8'd238:begin G_h <=4'd2;G_d<=4'd3;G_u<=4'd8;end
8'd239:begin G_h <=4'd2;G_d<=4'd3;G_u<=4'd9;end
8'd240:begin G_h <=4'd2;G_d<=4'd4;G_u<=4'd0;end
8'd241:begin G_h <=4'd2;G_d<=4'd4;G_u<=4'd1;end
8'd242:begin G_h <=4'd2;G_d<=4'd4;G_u<=4'd2;end
8'd243:begin G_h <=4'd2;G_d<=4'd4;G_u<=4'd3;end
8'd244:begin G_h <=4'd2;G_d<=4'd4;G_u<=4'd4;end
8'd245:begin G_h <=4'd2;G_d<=4'd4;G_u<=4'd5;end
8'd246:begin G_h <=4'd2;G_d<=4'd4;G_u<=4'd6;end
8'd247:begin G_h <=4'd2;G_d<=4'd4;G_u<=4'd7;end
8'd248:begin G_h <=4'd2;G_d<=4'd4;G_u<=4'd8;end
8'd249:begin G_h <=4'd2;G_d<=4'd4;G_u<=4'd9;end
8'd250:begin G_h <=4'd2;G_d<=4'd5;G_u<=4'd0;end
8'd251:begin G_h <=4'd2;G_d<=4'd5;G_u<=4'd1;end
8'd252:begin G_h <=4'd2;G_d<=4'd5;G_u<=4'd2;end
8'd253:begin G_h <=4'd2;G_d<=4'd5;G_u<=4'd3;end
8'd254:begin G_h <=4'd2;G_d<=4'd5;G_u<=4'd4;end
8'd255:begin G_h <=4'd2;G_d<=4'd5;G_u<=4'd5;end
endcase
end
always@(*)begin
case (B_detect)
8'd0:begin B_h <=4'd0;B_d<=4'd0;B_u<=4'd0;end
8'd1:begin B_h <=4'd0;B_d<=4'd0;B_u<=4'd1;end
8'd2:begin B_h <=4'd0;B_d<=4'd0;B_u<=4'd2;end
8'd3:begin B_h <=4'd0;B_d<=4'd0;B_u<=4'd3;end
8'd4:begin B_h <=4'd0;B_d<=4'd0;B_u<=4'd4;end
8'd5:begin B_h <=4'd0;B_d<=4'd0;B_u<=4'd5;end
8'd6:begin B_h <=4'd0;B_d<=4'd0;B_u<=4'd6;end
8'd7:begin B_h <=4'd0;B_d<=4'd0;B_u<=4'd7;end
8'd8:begin B_h <=4'd0;B_d<=4'd0;B_u<=4'd8;end
8'd9:begin B_h <=4'd0;B_d<=4'd0;B_u<=4'd9;end
8'd10:begin B_h <=4'd0;B_d<=4'd1;B_u<=4'd0;end
8'd11:begin B_h <=4'd0;B_d<=4'd1;B_u<=4'd1;end
8'd12:begin B_h <=4'd0;B_d<=4'd1;B_u<=4'd2;end
8'd13:begin B_h <=4'd0;B_d<=4'd1;B_u<=4'd3;end
8'd14:begin B_h <=4'd0;B_d<=4'd1;B_u<=4'd4;end
8'd15:begin B_h <=4'd0;B_d<=4'd1;B_u<=4'd5;end
8'd16:begin B_h <=4'd0;B_d<=4'd1;B_u<=4'd6;end
8'd17:begin B_h <=4'd0;B_d<=4'd1;B_u<=4'd7;end
8'd18:begin B_h <=4'd0;B_d<=4'd1;B_u<=4'd8;end
8'd19:begin B_h <=4'd0;B_d<=4'd1;B_u<=4'd9;end
8'd20:begin B_h <=4'd0;B_d<=4'd2;B_u<=4'd0;end
8'd21:begin B_h <=4'd0;B_d<=4'd2;B_u<=4'd1;end
8'd22:begin B_h <=4'd0;B_d<=4'd2;B_u<=4'd2;end
8'd23:begin B_h <=4'd0;B_d<=4'd2;B_u<=4'd3;end
8'd24:begin B_h <=4'd0;B_d<=4'd2;B_u<=4'd4;end
8'd25:begin B_h <=4'd0;B_d<=4'd2;B_u<=4'd5;end
8'd26:begin B_h <=4'd0;B_d<=4'd2;B_u<=4'd6;end
8'd27:begin B_h <=4'd0;B_d<=4'd2;B_u<=4'd7;end
8'd28:begin B_h <=4'd0;B_d<=4'd2;B_u<=4'd8;end
8'd29:begin B_h <=4'd0;B_d<=4'd2;B_u<=4'd9;end
8'd30:begin B_h <=4'd0;B_d<=4'd3;B_u<=4'd0;end
8'd31:begin B_h <=4'd0;B_d<=4'd3;B_u<=4'd1;end
8'd32:begin B_h <=4'd0;B_d<=4'd3;B_u<=4'd2;end
8'd33:begin B_h <=4'd0;B_d<=4'd3;B_u<=4'd3;end
8'd34:begin B_h <=4'd0;B_d<=4'd3;B_u<=4'd4;end
8'd35:begin B_h <=4'd0;B_d<=4'd3;B_u<=4'd5;end
8'd36:begin B_h <=4'd0;B_d<=4'd3;B_u<=4'd6;end
8'd37:begin B_h <=4'd0;B_d<=4'd3;B_u<=4'd7;end
8'd38:begin B_h <=4'd0;B_d<=4'd3;B_u<=4'd8;end
8'd39:begin B_h <=4'd0;B_d<=4'd3;B_u<=4'd9;end
8'd40:begin B_h <=4'd0;B_d<=4'd4;B_u<=4'd0;end
8'd41:begin B_h <=4'd0;B_d<=4'd4;B_u<=4'd1;end
8'd42:begin B_h <=4'd0;B_d<=4'd4;B_u<=4'd2;end
8'd43:begin B_h <=4'd0;B_d<=4'd4;B_u<=4'd3;end
8'd44:begin B_h <=4'd0;B_d<=4'd4;B_u<=4'd4;end
8'd45:begin B_h <=4'd0;B_d<=4'd4;B_u<=4'd5;end
8'd46:begin B_h <=4'd0;B_d<=4'd4;B_u<=4'd6;end
8'd47:begin B_h <=4'd0;B_d<=4'd4;B_u<=4'd7;end
8'd48:begin B_h <=4'd0;B_d<=4'd4;B_u<=4'd8;end
8'd49:begin B_h <=4'd0;B_d<=4'd4;B_u<=4'd9;end
8'd50:begin B_h <=4'd0;B_d<=4'd5;B_u<=4'd0;end
8'd51:begin B_h <=4'd0;B_d<=4'd5;B_u<=4'd1;end
8'd52:begin B_h <=4'd0;B_d<=4'd5;B_u<=4'd2;end
8'd53:begin B_h <=4'd0;B_d<=4'd5;B_u<=4'd3;end
8'd54:begin B_h <=4'd0;B_d<=4'd5;B_u<=4'd4;end
8'd55:begin B_h <=4'd0;B_d<=4'd5;B_u<=4'd5;end
8'd56:begin B_h <=4'd0;B_d<=4'd5;B_u<=4'd6;end
8'd57:begin B_h <=4'd0;B_d<=4'd5;B_u<=4'd7;end
8'd58:begin B_h <=4'd0;B_d<=4'd5;B_u<=4'd8;end
8'd59:begin B_h <=4'd0;B_d<=4'd5;B_u<=4'd9;end
8'd60:begin B_h <=4'd0;B_d<=4'd6;B_u<=4'd0;end
8'd61:begin B_h <=4'd0;B_d<=4'd6;B_u<=4'd1;end
8'd62:begin B_h <=4'd0;B_d<=4'd6;B_u<=4'd2;end
8'd63:begin B_h <=4'd0;B_d<=4'd6;B_u<=4'd3;end
8'd64:begin B_h <=4'd0;B_d<=4'd6;B_u<=4'd4;end
8'd65:begin B_h <=4'd0;B_d<=4'd6;B_u<=4'd5;end
8'd66:begin B_h <=4'd0;B_d<=4'd6;B_u<=4'd6;end
8'd67:begin B_h <=4'd0;B_d<=4'd6;B_u<=4'd7;end
8'd68:begin B_h <=4'd0;B_d<=4'd6;B_u<=4'd8;end
8'd69:begin B_h <=4'd0;B_d<=4'd6;B_u<=4'd9;end
8'd70:begin B_h <=4'd0;B_d<=4'd7;B_u<=4'd0;end
8'd71:begin B_h <=4'd0;B_d<=4'd7;B_u<=4'd1;end
8'd72:begin B_h <=4'd0;B_d<=4'd7;B_u<=4'd2;end
8'd73:begin B_h <=4'd0;B_d<=4'd7;B_u<=4'd3;end
8'd74:begin B_h <=4'd0;B_d<=4'd7;B_u<=4'd4;end
8'd75:begin B_h <=4'd0;B_d<=4'd7;B_u<=4'd5;end
8'd76:begin B_h <=4'd0;B_d<=4'd7;B_u<=4'd6;end
8'd77:begin B_h <=4'd0;B_d<=4'd7;B_u<=4'd7;end
8'd78:begin B_h <=4'd0;B_d<=4'd7;B_u<=4'd8;end
8'd79:begin B_h <=4'd0;B_d<=4'd7;B_u<=4'd9;end
8'd80:begin B_h <=4'd0;B_d<=4'd8;B_u<=4'd0;end
8'd81:begin B_h <=4'd0;B_d<=4'd8;B_u<=4'd1;end
8'd82:begin B_h <=4'd0;B_d<=4'd8;B_u<=4'd2;end
8'd83:begin B_h <=4'd0;B_d<=4'd8;B_u<=4'd3;end
8'd84:begin B_h <=4'd0;B_d<=4'd8;B_u<=4'd4;end
8'd85:begin B_h <=4'd0;B_d<=4'd8;B_u<=4'd5;end
8'd86:begin B_h <=4'd0;B_d<=4'd8;B_u<=4'd6;end
8'd87:begin B_h <=4'd0;B_d<=4'd8;B_u<=4'd7;end
8'd88:begin B_h <=4'd0;B_d<=4'd8;B_u<=4'd8;end
8'd89:begin B_h <=4'd0;B_d<=4'd8;B_u<=4'd9;end
8'd90:begin B_h <=4'd0;B_d<=4'd9;B_u<=4'd0;end
8'd91:begin B_h <=4'd0;B_d<=4'd9;B_u<=4'd1;end
8'd92:begin B_h <=4'd0;B_d<=4'd9;B_u<=4'd2;end
8'd93:begin B_h <=4'd0;B_d<=4'd9;B_u<=4'd3;end
8'd94:begin B_h <=4'd0;B_d<=4'd9;B_u<=4'd4;end
8'd95:begin B_h <=4'd0;B_d<=4'd9;B_u<=4'd5;end
8'd96:begin B_h <=4'd0;B_d<=4'd9;B_u<=4'd6;end
8'd97:begin B_h <=4'd0;B_d<=4'd9;B_u<=4'd7;end
8'd98:begin B_h <=4'd0;B_d<=4'd9;B_u<=4'd8;end
8'd99:begin B_h <=4'd0;B_d<=4'd9;B_u<=4'd9;end
8'd100:begin B_h <=4'd1;B_d<=4'd0;B_u<=4'd0;end
8'd101:begin B_h <=4'd1;B_d<=4'd0;B_u<=4'd1;end
8'd102:begin B_h <=4'd1;B_d<=4'd0;B_u<=4'd2;end
8'd103:begin B_h <=4'd1;B_d<=4'd0;B_u<=4'd3;end
8'd104:begin B_h <=4'd1;B_d<=4'd0;B_u<=4'd4;end
8'd105:begin B_h <=4'd1;B_d<=4'd0;B_u<=4'd5;end
8'd106:begin B_h <=4'd1;B_d<=4'd0;B_u<=4'd6;end
8'd107:begin B_h <=4'd1;B_d<=4'd0;B_u<=4'd7;end
8'd108:begin B_h <=4'd1;B_d<=4'd0;B_u<=4'd8;end
8'd109:begin B_h <=4'd1;B_d<=4'd0;B_u<=4'd9;end
8'd110:begin B_h <=4'd1;B_d<=4'd1;B_u<=4'd0;end
8'd111:begin B_h <=4'd1;B_d<=4'd1;B_u<=4'd1;end
8'd112:begin B_h <=4'd1;B_d<=4'd1;B_u<=4'd2;end
8'd113:begin B_h <=4'd1;B_d<=4'd1;B_u<=4'd3;end
8'd114:begin B_h <=4'd1;B_d<=4'd1;B_u<=4'd4;end
8'd115:begin B_h <=4'd1;B_d<=4'd1;B_u<=4'd5;end
8'd116:begin B_h <=4'd1;B_d<=4'd1;B_u<=4'd6;end
8'd117:begin B_h <=4'd1;B_d<=4'd1;B_u<=4'd7;end
8'd118:begin B_h <=4'd1;B_d<=4'd1;B_u<=4'd8;end
8'd119:begin B_h <=4'd1;B_d<=4'd1;B_u<=4'd9;end
8'd120:begin B_h <=4'd1;B_d<=4'd2;B_u<=4'd0;end
8'd121:begin B_h <=4'd1;B_d<=4'd2;B_u<=4'd1;end
8'd122:begin B_h <=4'd1;B_d<=4'd2;B_u<=4'd2;end
8'd123:begin B_h <=4'd1;B_d<=4'd2;B_u<=4'd3;end
8'd124:begin B_h <=4'd1;B_d<=4'd2;B_u<=4'd4;end
8'd125:begin B_h <=4'd1;B_d<=4'd2;B_u<=4'd5;end
8'd126:begin B_h <=4'd1;B_d<=4'd2;B_u<=4'd6;end
8'd127:begin B_h <=4'd1;B_d<=4'd2;B_u<=4'd7;end
8'd128:begin B_h <=4'd1;B_d<=4'd2;B_u<=4'd8;end
8'd129:begin B_h <=4'd1;B_d<=4'd2;B_u<=4'd9;end
8'd130:begin B_h <=4'd1;B_d<=4'd3;B_u<=4'd0;end
8'd131:begin B_h <=4'd1;B_d<=4'd3;B_u<=4'd1;end
8'd132:begin B_h <=4'd1;B_d<=4'd3;B_u<=4'd2;end
8'd133:begin B_h <=4'd1;B_d<=4'd3;B_u<=4'd3;end
8'd134:begin B_h <=4'd1;B_d<=4'd3;B_u<=4'd4;end
8'd135:begin B_h <=4'd1;B_d<=4'd3;B_u<=4'd5;end
8'd136:begin B_h <=4'd1;B_d<=4'd3;B_u<=4'd6;end
8'd137:begin B_h <=4'd1;B_d<=4'd3;B_u<=4'd7;end
8'd138:begin B_h <=4'd1;B_d<=4'd3;B_u<=4'd8;end
8'd139:begin B_h <=4'd1;B_d<=4'd3;B_u<=4'd9;end
8'd140:begin B_h <=4'd1;B_d<=4'd4;B_u<=4'd0;end
8'd141:begin B_h <=4'd1;B_d<=4'd4;B_u<=4'd1;end
8'd142:begin B_h <=4'd1;B_d<=4'd4;B_u<=4'd2;end
8'd143:begin B_h <=4'd1;B_d<=4'd4;B_u<=4'd3;end
8'd144:begin B_h <=4'd1;B_d<=4'd4;B_u<=4'd4;end
8'd145:begin B_h <=4'd1;B_d<=4'd4;B_u<=4'd5;end
8'd146:begin B_h <=4'd1;B_d<=4'd4;B_u<=4'd6;end
8'd147:begin B_h <=4'd1;B_d<=4'd4;B_u<=4'd7;end
8'd148:begin B_h <=4'd1;B_d<=4'd4;B_u<=4'd8;end
8'd149:begin B_h <=4'd1;B_d<=4'd4;B_u<=4'd9;end
8'd150:begin B_h <=4'd1;B_d<=4'd5;B_u<=4'd0;end
8'd151:begin B_h <=4'd1;B_d<=4'd5;B_u<=4'd1;end
8'd152:begin B_h <=4'd1;B_d<=4'd5;B_u<=4'd2;end
8'd153:begin B_h <=4'd1;B_d<=4'd5;B_u<=4'd3;end
8'd154:begin B_h <=4'd1;B_d<=4'd5;B_u<=4'd4;end
8'd155:begin B_h <=4'd1;B_d<=4'd5;B_u<=4'd5;end
8'd156:begin B_h <=4'd1;B_d<=4'd5;B_u<=4'd6;end
8'd157:begin B_h <=4'd1;B_d<=4'd5;B_u<=4'd7;end
8'd158:begin B_h <=4'd1;B_d<=4'd5;B_u<=4'd8;end
8'd159:begin B_h <=4'd1;B_d<=4'd5;B_u<=4'd9;end
8'd160:begin B_h <=4'd1;B_d<=4'd6;B_u<=4'd0;end
8'd161:begin B_h <=4'd1;B_d<=4'd6;B_u<=4'd1;end
8'd162:begin B_h <=4'd1;B_d<=4'd6;B_u<=4'd2;end
8'd163:begin B_h <=4'd1;B_d<=4'd6;B_u<=4'd3;end
8'd164:begin B_h <=4'd1;B_d<=4'd6;B_u<=4'd4;end
8'd165:begin B_h <=4'd1;B_d<=4'd6;B_u<=4'd5;end
8'd166:begin B_h <=4'd1;B_d<=4'd6;B_u<=4'd6;end
8'd167:begin B_h <=4'd1;B_d<=4'd6;B_u<=4'd7;end
8'd168:begin B_h <=4'd1;B_d<=4'd6;B_u<=4'd8;end
8'd169:begin B_h <=4'd1;B_d<=4'd6;B_u<=4'd9;end
8'd170:begin B_h <=4'd1;B_d<=4'd7;B_u<=4'd0;end
8'd171:begin B_h <=4'd1;B_d<=4'd7;B_u<=4'd1;end
8'd172:begin B_h <=4'd1;B_d<=4'd7;B_u<=4'd2;end
8'd173:begin B_h <=4'd1;B_d<=4'd7;B_u<=4'd3;end
8'd174:begin B_h <=4'd1;B_d<=4'd7;B_u<=4'd4;end
8'd175:begin B_h <=4'd1;B_d<=4'd7;B_u<=4'd5;end
8'd176:begin B_h <=4'd1;B_d<=4'd7;B_u<=4'd6;end
8'd177:begin B_h <=4'd1;B_d<=4'd7;B_u<=4'd7;end
8'd178:begin B_h <=4'd1;B_d<=4'd7;B_u<=4'd8;end
8'd179:begin B_h <=4'd1;B_d<=4'd7;B_u<=4'd9;end
8'd180:begin B_h <=4'd1;B_d<=4'd8;B_u<=4'd0;end
8'd181:begin B_h <=4'd1;B_d<=4'd8;B_u<=4'd1;end
8'd182:begin B_h <=4'd1;B_d<=4'd8;B_u<=4'd2;end
8'd183:begin B_h <=4'd1;B_d<=4'd8;B_u<=4'd3;end
8'd184:begin B_h <=4'd1;B_d<=4'd8;B_u<=4'd4;end
8'd185:begin B_h <=4'd1;B_d<=4'd8;B_u<=4'd5;end
8'd186:begin B_h <=4'd1;B_d<=4'd8;B_u<=4'd6;end
8'd187:begin B_h <=4'd1;B_d<=4'd8;B_u<=4'd7;end
8'd188:begin B_h <=4'd1;B_d<=4'd8;B_u<=4'd8;end
8'd189:begin B_h <=4'd1;B_d<=4'd8;B_u<=4'd9;end
8'd190:begin B_h <=4'd1;B_d<=4'd9;B_u<=4'd0;end
8'd191:begin B_h <=4'd1;B_d<=4'd9;B_u<=4'd1;end
8'd192:begin B_h <=4'd1;B_d<=4'd9;B_u<=4'd2;end
8'd193:begin B_h <=4'd1;B_d<=4'd9;B_u<=4'd3;end
8'd194:begin B_h <=4'd1;B_d<=4'd9;B_u<=4'd4;end
8'd195:begin B_h <=4'd1;B_d<=4'd9;B_u<=4'd5;end
8'd196:begin B_h <=4'd1;B_d<=4'd9;B_u<=4'd6;end
8'd197:begin B_h <=4'd1;B_d<=4'd9;B_u<=4'd7;end
8'd198:begin B_h <=4'd1;B_d<=4'd9;B_u<=4'd8;end
8'd199:begin B_h <=4'd1;B_d<=4'd9;B_u<=4'd9;end
8'd200:begin B_h <=4'd2;B_d<=4'd0;B_u<=4'd0;end
8'd201:begin B_h <=4'd2;B_d<=4'd0;B_u<=4'd1;end
8'd202:begin B_h <=4'd2;B_d<=4'd0;B_u<=4'd2;end
8'd203:begin B_h <=4'd2;B_d<=4'd0;B_u<=4'd3;end
8'd204:begin B_h <=4'd2;B_d<=4'd0;B_u<=4'd4;end
8'd205:begin B_h <=4'd2;B_d<=4'd0;B_u<=4'd5;end
8'd206:begin B_h <=4'd2;B_d<=4'd0;B_u<=4'd6;end
8'd207:begin B_h <=4'd2;B_d<=4'd0;B_u<=4'd7;end
8'd208:begin B_h <=4'd2;B_d<=4'd0;B_u<=4'd8;end
8'd209:begin B_h <=4'd2;B_d<=4'd0;B_u<=4'd9;end
8'd210:begin B_h <=4'd2;B_d<=4'd1;B_u<=4'd0;end
8'd211:begin B_h <=4'd2;B_d<=4'd1;B_u<=4'd1;end
8'd212:begin B_h <=4'd2;B_d<=4'd1;B_u<=4'd2;end
8'd213:begin B_h <=4'd2;B_d<=4'd1;B_u<=4'd3;end
8'd214:begin B_h <=4'd2;B_d<=4'd1;B_u<=4'd4;end
8'd215:begin B_h <=4'd2;B_d<=4'd1;B_u<=4'd5;end
8'd216:begin B_h <=4'd2;B_d<=4'd1;B_u<=4'd6;end
8'd217:begin B_h <=4'd2;B_d<=4'd1;B_u<=4'd7;end
8'd218:begin B_h <=4'd2;B_d<=4'd1;B_u<=4'd8;end
8'd219:begin B_h <=4'd2;B_d<=4'd1;B_u<=4'd9;end
8'd220:begin B_h <=4'd2;B_d<=4'd2;B_u<=4'd0;end
8'd221:begin B_h <=4'd2;B_d<=4'd2;B_u<=4'd1;end
8'd222:begin B_h <=4'd2;B_d<=4'd2;B_u<=4'd2;end
8'd223:begin B_h <=4'd2;B_d<=4'd2;B_u<=4'd3;end
8'd224:begin B_h <=4'd2;B_d<=4'd2;B_u<=4'd4;end
8'd225:begin B_h <=4'd2;B_d<=4'd2;B_u<=4'd5;end
8'd226:begin B_h <=4'd2;B_d<=4'd2;B_u<=4'd6;end
8'd227:begin B_h <=4'd2;B_d<=4'd2;B_u<=4'd7;end
8'd228:begin B_h <=4'd2;B_d<=4'd2;B_u<=4'd8;end
8'd229:begin B_h <=4'd2;B_d<=4'd2;B_u<=4'd9;end
8'd230:begin B_h <=4'd2;B_d<=4'd3;B_u<=4'd0;end
8'd231:begin B_h <=4'd2;B_d<=4'd3;B_u<=4'd1;end
8'd232:begin B_h <=4'd2;B_d<=4'd3;B_u<=4'd2;end
8'd233:begin B_h <=4'd2;B_d<=4'd3;B_u<=4'd3;end
8'd234:begin B_h <=4'd2;B_d<=4'd3;B_u<=4'd4;end
8'd235:begin B_h <=4'd2;B_d<=4'd3;B_u<=4'd5;end
8'd236:begin B_h <=4'd2;B_d<=4'd3;B_u<=4'd6;end
8'd237:begin B_h <=4'd2;B_d<=4'd3;B_u<=4'd7;end
8'd238:begin B_h <=4'd2;B_d<=4'd3;B_u<=4'd8;end
8'd239:begin B_h <=4'd2;B_d<=4'd3;B_u<=4'd9;end
8'd240:begin B_h <=4'd2;B_d<=4'd4;B_u<=4'd0;end
8'd241:begin B_h <=4'd2;B_d<=4'd4;B_u<=4'd1;end
8'd242:begin B_h <=4'd2;B_d<=4'd4;B_u<=4'd2;end
8'd243:begin B_h <=4'd2;B_d<=4'd4;B_u<=4'd3;end
8'd244:begin B_h <=4'd2;B_d<=4'd4;B_u<=4'd4;end
8'd245:begin B_h <=4'd2;B_d<=4'd4;B_u<=4'd5;end
8'd246:begin B_h <=4'd2;B_d<=4'd4;B_u<=4'd6;end
8'd247:begin B_h <=4'd2;B_d<=4'd4;B_u<=4'd7;end
8'd248:begin B_h <=4'd2;B_d<=4'd4;B_u<=4'd8;end
8'd249:begin B_h <=4'd2;B_d<=4'd4;B_u<=4'd9;end
8'd250:begin B_h <=4'd2;B_d<=4'd5;B_u<=4'd0;end
8'd251:begin B_h <=4'd2;B_d<=4'd5;B_u<=4'd1;end
8'd252:begin B_h <=4'd2;B_d<=4'd5;B_u<=4'd2;end
8'd253:begin B_h <=4'd2;B_d<=4'd5;B_u<=4'd3;end
8'd254:begin B_h <=4'd2;B_d<=4'd5;B_u<=4'd4;end
8'd255:begin B_h <=4'd2;B_d<=4'd5;B_u<=4'd5;end
endcase
end
 
endmodule
